library verilog;
use verilog.vl_types.all;
entity tb_mbe_mult is
end tb_mbe_mult;
