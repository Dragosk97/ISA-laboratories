library verilog;
use verilog.vl_types.all;
entity tb_m is
end tb_m;
