library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity datapath is
    port ( 

    
    );
end datapath;

ARCHITECTURE structural of datapath is

begin

end structural;